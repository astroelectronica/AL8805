.title KiCad schematic
.include "C:/AE/AL8805/_models/AL8805.spice.txt"
.include "C:/AE/AL8805/_models/C2012X5R1H475K125AB_p.mod"
.include "C:/AE/AL8805/_models/C2012X7R2A104K125AE_p.mod"
.include "C:/AE/AL8805/_models/C3225X7T2J104M160AC_p.mod"
.include "C:/AE/AL8805/_models/DFLS240L.spice.txt"
.include "C:/AE/AL8805/_models/TPC_1028_744065330_33u.lib"
.include "C:/AE/AL8805/_models/XPE_SPICE.lib"
D4 /LDB4 /LDB5 XLampXPEgreen
V2 VCC 0 {VSOURCE}
D2 /A /LDB3 XLampXPEgreen
D3 /LDB3 /LDB4 XLampXPEgreen
XU4 /A /K C3225X7T2J104M160AC_p
XU5 /K /SW TPC_1028_744065330_33u
D5 /LDB5 /LDB6 XLampXPEgreen
D6 /LDB6 /K XLampXPEgreen
R2 VCC /A {RSENSE2}
R1 VCC /A {RSENSE1}
XU1 /SW 0 /CTRL /A VCC AL8805
D1 /SW VCC DI_DFLS240L
V1 /PWM 0  PULSE(0 {VPUL} {DELAY} {TR} {TF} {DUTY} {CYCLE})
XU3 VCC 0 C2012X7R2A104K125AE_p
R3 /PWM /CTRL {RCTRL}
XU2 VCC 0 C2012X5R1H475K125AB_p
.end
